module with_parameter_port_list #(
        P1,
        localparam L2 = P1+1,
        parameter P2)
        ( /*port list...*/ );
        parameter  L3 = "synonym for the localparam";
        localparam L4 = "localparam";
        // ...
endmodule