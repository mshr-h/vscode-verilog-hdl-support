module float_add (
);

endmodule

module test (
);
float_add fa (
);

endmodule
