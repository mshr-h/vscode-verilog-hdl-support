module test (
);

endmodulea

module float_add (
);

endmodule

// % iverilog -t null 01_sntax_error.v                                     
// 01_sntax_error.yv:6: syntax error
// 01_syntax_error.v:4: error: Invalid module instantiation
